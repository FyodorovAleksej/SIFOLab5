lpm_constant8_inst : lpm_constant8 PORT MAP (
		result	 => result_sig
	);
