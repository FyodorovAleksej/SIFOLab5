lpm_constant11_inst : lpm_constant11 PORT MAP (
		result	 => result_sig
	);
