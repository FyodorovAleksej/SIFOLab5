lpm_constant7_inst : lpm_constant7 PORT MAP (
		result	 => result_sig
	);
