lpm_constant6_inst : lpm_constant6 PORT MAP (
		result	 => result_sig
	);
