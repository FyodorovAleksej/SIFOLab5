lpm_compare0_inst : lpm_compare0 PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		AeB	 => AeB_sig
	);
