lpm_or0_inst : lpm_or0 PORT MAP (
		data0x	 => data0x_sig,
		data1x	 => data1x_sig,
		result	 => result_sig
	);
