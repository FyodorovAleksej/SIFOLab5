lpm_constant9_inst : lpm_constant9 PORT MAP (
		result	 => result_sig
	);
