lpm_constant1_inst : lpm_constant1 PORT MAP (
		result	 => result_sig
	);
