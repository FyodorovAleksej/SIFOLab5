lpm_constant4_inst : lpm_constant4 PORT MAP (
		result	 => result_sig
	);
