lpm_constant5_inst : lpm_constant5 PORT MAP (
		result	 => result_sig
	);
