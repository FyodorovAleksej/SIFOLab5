lpm_constant10_inst : lpm_constant10 PORT MAP (
		result	 => result_sig
	);
